(* dont_touch = "true" *)

import control_pkg::*;

`timescale 1ns/1ps

module aludec (
    
    input logic         opb5, // for sub detection
    input logic  [2:0]  funct3,
    input logic         funct7b5, // instr[30] for SUB/SRA
    input logic  [1:0]  ALUOp,
    output logic [3:0]  ALUControl
    
);

    logic RtypeSub;
    assign RtypeSub = funct7b5 & opb5; // TRUE for R-type SUB

    always_comb begin

        unique case (ALUOp)

            2'b00: begin

                ALUControl = ADD; // load/store, addi
                    
            end

            2'b01: begin

                ALUControl = SUB; // branches
                    
            end

            default: begin

                unique case (funct3)
                    
                    3'b000: ALUControl = RtypeSub ? SUB : ADD; // same for rv32 & rv64
                    3'b001: ALUControl = SLL; // same for rv32 & rv64
                    3'b010: ALUControl = SLT; // slt/slti (signed)
                    3'b011: ALUControl = SLTU; // sltu/sltiu (unsigned)
                    3'b100: ALUControl = XOR;
                    3'b101: ALUControl = funct7b5 ? SRA : SRL; // sra/srai or srl/srli (same for rv32 & rv64)
                    3'b110: ALUControl = OR; // or/ori
                    3'b111: ALUControl = AND; // and/andi

                endcase

            end

        endcase

    end

endmodule